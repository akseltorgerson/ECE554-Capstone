module proc();


endmodule