module fetch_stage(clk, rst, halt, insr, pcplus4, next_pc);

endmodule