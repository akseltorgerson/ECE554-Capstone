module twiddle_ROM();
    
endmodule