module fft_accel(
    input clk, rst, startF, startI, loadF, filter,
    input [17:0] sigNum,
    output done, calculating
);

    ////////////////////////
    ////// modules//////////
    ////////////////////////
    twiddle_ROM rom1()


endmodule